Linear DWDM Link
Ra 1 2 NODE_ADD NLOSS=14.0
Ab 2 3 EDFA_BOOSTER
L1 3 4 OPTLINK_NZ LEN=40.0
R1 4 5 NODE2 NLOSS=16.0
L2 5 6 OPTLINK_NZ LEN=40.0
Ap 6 7 EDFA_PRE
Rd 7 8 NODE_DROP NLOSS=15.0

Pin 1 0 0
.optqpt

.MODEL OPTLINK_SM L(ALPHA=0.27 D=-17.0)
.MODEL OPTLINK_NZ L(ALPHA=0.22 D=-10.0)
.MODEL EDFA_BOOSTER A(G=23 NF=5.5 LOSS =1)
.MODEL EDFA_LINE A(G=20 NF=5 LOSS =1)
.MODEL EDFA_PRE A(G=20 NF=6 LOSS =1)
.MODEL NODE_ADD R(NLOSS=14.0)
.MODEL NODE1 R(NLOSS=14)
.MODEL NODE2 R(NLOSS=16)
.MODEL NODE3 R(NLOSS=18)
.MODEL NODE_DROP R(NLOSS=15.0)
.MODEL DISP_30Km D(PL=4 DC=510)
.MODEL DISP_60Km D(PL=4 DC=1020)
.MODEL DISP_80Km D(PL=4 DC=1360)
.MODEL DISP_120Km D(PL=4 DC=2040)


.end