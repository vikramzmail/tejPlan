Linear DWDM Link
L1 1 2 OPTLINK LEN=125
A1 2 3 EDFA
L2 3 4 OPTLINK LEN=125
A2 4 5 EDFA
L3 5 6 OPTLINK LEN=125
A3 6 7 EDFA
L4 7 8 OPTLINK LEN=125

Pin 1 0 0
.optqpt

.MODEL OPTLINK L(ALPHA=0.2 D=-17.0)
.MODEL EDFA A(G=22 NF=5 LOSS =1)


.end